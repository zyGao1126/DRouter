VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
 DATABASE MICRONS 2000 ;
END UNITS

LAYER TEXT
 TYPE MASTERSLICE ;
END TEXT

LAYER METAL1
 TYPE ROUTING ;
 PITCH 0.41 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.16 ;
 MINWIDTH 0.16 ;
 SPACING 0.18 ;
END METAL1

LAYER VIA12
 TYPE CUT ;
 SPACING 0.22 ;
END VIA12

LAYER METAL2
 TYPE ROUTING ;
 PITCH 0.46 ;
 DIRECTION VERTICAL ;
 WIDTH 0.2 ;
 MINWIDTH 0.2 ;
 SPACING 0.21 ;
 AREA 0.144 ;
END METAL2

LAYER VIA23
 TYPE CUT ;
 SPACING 0.22 ;
END VIA23

LAYER METAL3
 TYPE ROUTING ;
 PITCH 0.41 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.2 ;
 MINWIDTH 0.2 ;
 SPACING 0.21 ;
 AREA 0.144 ;
END METAL3

LAYER VIA34
 TYPE CUT ;
 SPACING 0.22 ;
END VIA34

LAYER METAL4
 TYPE ROUTING ;
 PITCH 0.46 ;
 DIRECTION VERTICAL ;
 WIDTH 0.2 ;
 MINWIDTH 0.2 ;
 SPACING 0.21 ;
 AREA 0.144 ;
END METAL4

LAYER VIA45
 TYPE CUT ;
 SPACING 0.22 ;
END VIA45

LAYER METAL5
 TYPE ROUTING ;
 PITCH 0.41 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.2 ;
 MINWIDTH 0.2 ;
 SPACING 0.21 ;
 AREA 0.144 ;
END METAL5

LAYER VIA56
 TYPE CUT ;
 SPACING 0.22 ;
END VIA56

LAYER METAL6
 TYPE ROUTING ;
 PITCH 0.46 ;
 DIRECTION VERTICAL ;
 WIDTH 0.2 ;
 MINWIDTH 0.2 ;
 SPACING 0.21 ;
 AREA 0.144 ;
END METAL6

LAYER VIA67
 TYPE CUT ;
 SPACING 0.22 ;
END VIA67

LAYER METAL7
 TYPE ROUTING ;
 PITCH 0.41 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.2 ;
 MINWIDTH 0.2 ;
 SPACING 0.21 ; 
END METAL7

LAYER VIA78
 TYPE CUT ;
 SPACING 0.35 ;
END VIA78

LAYER METAL8
 TYPE ROUTING ;
 PITCH 1.38 ;
 DIRECTION VERTICAL ;
 WIDTH 0.44 ;
 MINWIDTH 0.44 ;
 SPACING 0.46 ;
END METAL8

VIARULE via1Array GENERATE
  LAYER METAL1 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER METAL2 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER VIA12 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END via1Array

VIARULE via2Array GENERATE
  LAYER METAL2 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER METAL3 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER VIA23 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END via2Array

VIARULE via3Array GENERATE
  LAYER METAL3 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER METAL4 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER VIA34 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END via3Array

VIARULE via4Array GENERATE
  LAYER METAL4 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER METAL5 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER VIA45 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END via4Array

VIARULE via5Array GENERATE
  LAYER METAL5 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER METAL6 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER VIA56 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END via5Array

VIARULE via6Array GENERATE
  LAYER METAL6 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER METAL7 ;
    ENCLOSURE 0.05 0.05 ;
  LAYER VIA67 ;
    RECT -0.095 -0.095 0.095 0.095 ;
    SPACING 0.48 BY 0.48 ;
END via6Array

VIARULE via7Array GENERATE
  LAYER METAL7 ;
    ENCLOSURE 0.05 0.09 ;
  LAYER METAL8 ;
    ENCLOSURE 0.05 0.09 ;
  LAYER VIA78 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.9 BY 0.9 ;
END via7Array

VIA via1 DEFAULT
  LAYER VIA12 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL1 ;
    RECT -0.105 -0.145 0.105 0.145 ;
  LAYER METAL2 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  END via1

VIA via1vh DEFAULT
  LAYER VIA12 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL1 ;
    RECT -0.105 -0.145 0.105 0.145 ;
  LAYER METAL2 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via1vh

VIA via2 DEFAULT
  LAYER VIA23 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL2 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  LAYER METAL3 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via2

VIA via2hh DEFAULT
  LAYER VIA23 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL2 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  LAYER METAL3 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via2hh

VIA via2ts DEFAULT
  LAYER VIA23 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL2 ;
    RECT -0.1 -0.36 0.1 0.36 ;
  LAYER METAL3 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via2ts

VIA via3 DEFAULT
  LAYER VIA34 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL3 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  LAYER METAL4 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  END via3

VIA via3hh DEFAULT
  LAYER VIA34 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL3 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  LAYER METAL4 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via3hh

VIA via3ts DEFAULT
  LAYER VIA34 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL3 ;
    RECT -0.36 -0.1 0.36 0.1 ;
  LAYER METAL4 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  END via3ts

VIA via4 DEFAULT
  LAYER VIA45 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL4 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  LAYER METAL5 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via4

VIA via4hh DEFAULT
  LAYER VIA45 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL4 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  LAYER METAL5 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via4hh

VIA via4ts DEFAULT
  LAYER VIA45 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL4 ;
    RECT -0.1 -0.36 0.1 0.36 ;
  LAYER METAL5 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via4ts

VIA via5 DEFAULT
  LAYER VIA56 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL5 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  LAYER METAL6 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  END via5

VIA via5vv DEFAULT
  LAYER VIA56 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL5 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  LAYER METAL6 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  END via5vv

VIA via5ts DEFAULT
  LAYER VIA56 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL5 ;
    RECT -0.36 -0.1 0.36 0.1 ;
  LAYER METAL6 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  END via5ts

VIA via6 DEFAULT
  LAYER VIA67 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL6 ;
    RECT -0.1 -0.145 0.1 0.145 ;
  LAYER METAL7 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via6

VIA via6hh DEFAULT
  LAYER VIA67 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL6 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  LAYER METAL7 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via6hh

VIA via6ts DEFAULT
  LAYER VIA67 ;
    RECT -0.095 -0.095 0.095 0.095 ;
  LAYER METAL6 ;
    RECT -0.1 -0.36 0.1 0.36 ;
  LAYER METAL7 ;
    RECT -0.145 -0.1 0.145 0.1 ;
  END via6ts

VIA via7 DEFAULT
  LAYER VIA78 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER METAL7 ;
    RECT -0.23 -0.19 0.23 0.19 ;
  LAYER METAL8 ;
    RECT -0.27 -0.27 0.27 0.27 ;
  END via7

MACRO CELL1
 CLASS CORE ;
 FOREIGN CELL1 ;
 ORIGIN 0 0 ;
 SIZE 14.26 BY 3.69 ;
 SYMMETRY X Y  ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER METAL1 ;
 RECT 1.505 1.275 1.745 1.535 ;
 RECT 1.505 1.535 1.715 1.83 ;
 END
 END SE

 PIN ECK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER METAL1 ;
 RECT 8.605 2.585 13.995 2.65 ;
 RECT 9.625 2.65 9.885 3.115 ;
 RECT 8.605 2.65 8.865 3.115 ;
 RECT 13.64 2.65 13.99 3.115 ;
 RECT 11.625 2.65 11.925 2.995 ;
 RECT 10.645 2.65 10.915 2.995 ;
 RECT 8.605 2.335 14.135 2.585 ;
 RECT 8.605 2.045 13.995 2.335 ;
 RECT 11.665 2.995 11.925 3.115 ;
 RECT 10.645 2.995 10.905 3.115 ;
 RECT 12.965 1.305 13.795 1.925 ;
 RECT 8.53 0.705 14.13 1.305 ;
 RECT 12.965 1.925 13.995 2.045 ;
 RECT 12.685 2.65 12.945 3.115 ;
 END
 END ECK

 PIN E
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER METAL1 ;
 RECT 1.965 1.755 2.23 1.825 ;
 RECT 1.94 1.825 2.38 2.035 ;
 RECT 1.965 1.7 2.175 1.755 ;
 END
 END E

 PIN CK
 DIRECTION INPUT ;
 USE CLOCK ;
 PORT
 LAYER METAL1 ;
 RECT 0.125 1.765 0.37 2.045 ;
 RECT 0.125 1.575 0.345 1.765 ;
 RECT 0.125 2.045 0.345 2.145 ;
 END
 END CK

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER METAL1 ;
 RECT 0 -0.25 14.26 0.25 ;
 RECT 12.325 0.25 12.585 0.405 ;
 RECT 11.31 0.25 11.57 0.405 ;
 RECT 10.255 0.25 10.515 0.405 ;
 RECT 9.22 0.25 9.48 0.405 ;
 RECT 8.185 0.25 8.445 0.405 ;
 RECT 7.17 0.25 7.43 0.405 ;
 RECT 6.125 0.25 6.385 0.405 ;
 RECT 4.575 0.25 5.295 0.405 ;
 RECT 2.325 0.25 2.925 0.405 ;
 RECT 0.675 0.25 1.275 0.405 ;
 RECT 0.675 0.405 0.935 0.755 ;
 RECT 13.355 0.25 13.615 0.405 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER METAL1 ;
 RECT 0 3.44 14.26 3.94 ;
 RECT 12.175 2.895 12.435 3.44 ;
 RECT 11.155 2.895 11.415 3.44 ;
 RECT 10.135 2.895 10.395 3.44 ;
 RECT 9.115 2.895 9.375 3.44 ;
 RECT 8.095 2.105 8.355 3.44 ;
 RECT 7.075 2.595 7.335 3.44 ;
 RECT 5.195 3.285 5.455 3.44 ;
 RECT 2.815 3.285 3.075 3.44 ;
 RECT 1.235 2.86 1.495 3.44 ;
 RECT 0.15 2.905 0.41 3.44 ;
 RECT 13.195 2.895 13.455 3.44 ;
 END
 END VDD

END CELL1

MACRO CELL2
 CLASS CORE ;
 FOREIGN CELL2 ;
 ORIGIN 0 0 ;
 SIZE 9.66 BY 3.69 ;
 SYMMETRY X Y  ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER METAL1 ;
 RECT 9.265 1.105 9.535 1.235 ;
 RECT 9.265 0.975 9.525 1.105 ;
 RECT 9.325 1.235 9.535 1.955 ;
 RECT 9.265 1.955 9.535 2.175 ;
 RECT 9.265 2.175 9.525 2.555 ;
 END
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER METAL1 ;
 RECT 1.64 1.29 2.175 1.55 ;
 RECT 1.965 1.55 2.175 1.58 ;
 END
 END D

 PIN CK
 DIRECTION INPUT ;
 USE CLOCK ;
 PORT
 LAYER METAL1 ;
 RECT 0.12 1.695 0.395 1.955 ;
 RECT 0.12 1.52 0.345 1.695 ;
 RECT 0.12 1.955 0.345 2.13 ;
 END
 END CK

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER METAL1 ;
 RECT 0 -0.25 9.66 0.25 ;
 RECT 7.565 0.25 7.825 1.045 ;
 RECT 5.625 0.25 5.885 0.405 ;
 RECT 4.375 0.25 4.635 0.405 ;
 RECT 2.475 0.25 2.635 0.745 ;
 RECT 0.705 0.25 1.305 0.405 ;
 RECT 8.755 0.25 9.015 1.235 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER METAL1 ;
 RECT 0 3.44 9.66 3.94 ;
 RECT 5.065 3.285 6.125 3.44 ;
 RECT 3.305 3.285 3.565 3.44 ;
 RECT 2.42 3.285 2.68 3.44 ;
 RECT 0.49 3.285 0.75 3.44 ;
 RECT 8.365 2.895 8.965 3.44 ;
 END
 END VDD

END CELL2

END LIBRARY
